`ifndef DATA_TYPE_SVH
`define DATA_TYPE_SVH

typedef struct packed {
  logic [3:0] value;
  logic       valid;      
} data_t;


`endif
