priority case(1'b1)
in[0] : out[0] = 1'b1;
in[1] : out[1] = 1'b1;
in[2] : out[2] = 1'b1;
in[3] : out[3] = 1'b1;
endcase
