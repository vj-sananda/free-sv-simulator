priority case(1'b1)
in[0] : out[0] = 1'b1;
in[1] : out[1] = 1'b1;
in[2] : out[2] = 1'b1;
in[3] : out[3] = 1'b1;
in[4] : out[4] = 1'b1;
in[5] : out[5] = 1'b1;
in[6] : out[6] = 1'b1;
in[7] : out[7] = 1'b1;
in[8] : out[8] = 1'b1;
in[9] : out[9] = 1'b1;
in[10] : out[10] = 1'b1;
in[11] : out[11] = 1'b1;
in[12] : out[12] = 1'b1;
in[13] : out[13] = 1'b1;
in[14] : out[14] = 1'b1;
in[15] : out[15] = 1'b1;
in[16] : out[16] = 1'b1;
in[17] : out[17] = 1'b1;
in[18] : out[18] = 1'b1;
in[19] : out[19] = 1'b1;
in[20] : out[20] = 1'b1;
in[21] : out[21] = 1'b1;
in[22] : out[22] = 1'b1;
in[23] : out[23] = 1'b1;
in[24] : out[24] = 1'b1;
in[25] : out[25] = 1'b1;
in[26] : out[26] = 1'b1;
in[27] : out[27] = 1'b1;
in[28] : out[28] = 1'b1;
in[29] : out[29] = 1'b1;
in[30] : out[30] = 1'b1;
in[31] : out[31] = 1'b1;
in[32] : out[32] = 1'b1;
in[33] : out[33] = 1'b1;
in[34] : out[34] = 1'b1;
in[35] : out[35] = 1'b1;
in[36] : out[36] = 1'b1;
in[37] : out[37] = 1'b1;
in[38] : out[38] = 1'b1;
in[39] : out[39] = 1'b1;
in[40] : out[40] = 1'b1;
in[41] : out[41] = 1'b1;
in[42] : out[42] = 1'b1;
in[43] : out[43] = 1'b1;
in[44] : out[44] = 1'b1;
in[45] : out[45] = 1'b1;
in[46] : out[46] = 1'b1;
in[47] : out[47] = 1'b1;
in[48] : out[48] = 1'b1;
in[49] : out[49] = 1'b1;
in[50] : out[50] = 1'b1;
in[51] : out[51] = 1'b1;
in[52] : out[52] = 1'b1;
in[53] : out[53] = 1'b1;
in[54] : out[54] = 1'b1;
in[55] : out[55] = 1'b1;
in[56] : out[56] = 1'b1;
in[57] : out[57] = 1'b1;
in[58] : out[58] = 1'b1;
in[59] : out[59] = 1'b1;
in[60] : out[60] = 1'b1;
in[61] : out[61] = 1'b1;
in[62] : out[62] = 1'b1;
in[63] : out[63] = 1'b1;
in[64] : out[64] = 1'b1;
in[65] : out[65] = 1'b1;
in[66] : out[66] = 1'b1;
in[67] : out[67] = 1'b1;
in[68] : out[68] = 1'b1;
in[69] : out[69] = 1'b1;
in[70] : out[70] = 1'b1;
in[71] : out[71] = 1'b1;
in[72] : out[72] = 1'b1;
in[73] : out[73] = 1'b1;
in[74] : out[74] = 1'b1;
in[75] : out[75] = 1'b1;
in[76] : out[76] = 1'b1;
in[77] : out[77] = 1'b1;
in[78] : out[78] = 1'b1;
in[79] : out[79] = 1'b1;
in[80] : out[80] = 1'b1;
in[81] : out[81] = 1'b1;
in[82] : out[82] = 1'b1;
in[83] : out[83] = 1'b1;
in[84] : out[84] = 1'b1;
in[85] : out[85] = 1'b1;
in[86] : out[86] = 1'b1;
in[87] : out[87] = 1'b1;
in[88] : out[88] = 1'b1;
in[89] : out[89] = 1'b1;
in[90] : out[90] = 1'b1;
in[91] : out[91] = 1'b1;
in[92] : out[92] = 1'b1;
in[93] : out[93] = 1'b1;
in[94] : out[94] = 1'b1;
in[95] : out[95] = 1'b1;
in[96] : out[96] = 1'b1;
in[97] : out[97] = 1'b1;
in[98] : out[98] = 1'b1;
in[99] : out[99] = 1'b1;
in[100] : out[100] = 1'b1;
in[101] : out[101] = 1'b1;
in[102] : out[102] = 1'b1;
in[103] : out[103] = 1'b1;
in[104] : out[104] = 1'b1;
in[105] : out[105] = 1'b1;
in[106] : out[106] = 1'b1;
in[107] : out[107] = 1'b1;
in[108] : out[108] = 1'b1;
in[109] : out[109] = 1'b1;
in[110] : out[110] = 1'b1;
in[111] : out[111] = 1'b1;
in[112] : out[112] = 1'b1;
in[113] : out[113] = 1'b1;
in[114] : out[114] = 1'b1;
in[115] : out[115] = 1'b1;
in[116] : out[116] = 1'b1;
in[117] : out[117] = 1'b1;
in[118] : out[118] = 1'b1;
in[119] : out[119] = 1'b1;
in[120] : out[120] = 1'b1;
in[121] : out[121] = 1'b1;
in[122] : out[122] = 1'b1;
in[123] : out[123] = 1'b1;
in[124] : out[124] = 1'b1;
in[125] : out[125] = 1'b1;
in[126] : out[126] = 1'b1;
in[127] : out[127] = 1'b1;
in[128] : out[128] = 1'b1;
in[129] : out[129] = 1'b1;
in[130] : out[130] = 1'b1;
in[131] : out[131] = 1'b1;
in[132] : out[132] = 1'b1;
in[133] : out[133] = 1'b1;
in[134] : out[134] = 1'b1;
in[135] : out[135] = 1'b1;
in[136] : out[136] = 1'b1;
in[137] : out[137] = 1'b1;
in[138] : out[138] = 1'b1;
in[139] : out[139] = 1'b1;
in[140] : out[140] = 1'b1;
in[141] : out[141] = 1'b1;
in[142] : out[142] = 1'b1;
in[143] : out[143] = 1'b1;
in[144] : out[144] = 1'b1;
in[145] : out[145] = 1'b1;
in[146] : out[146] = 1'b1;
in[147] : out[147] = 1'b1;
in[148] : out[148] = 1'b1;
in[149] : out[149] = 1'b1;
in[150] : out[150] = 1'b1;
in[151] : out[151] = 1'b1;
in[152] : out[152] = 1'b1;
in[153] : out[153] = 1'b1;
in[154] : out[154] = 1'b1;
in[155] : out[155] = 1'b1;
in[156] : out[156] = 1'b1;
in[157] : out[157] = 1'b1;
in[158] : out[158] = 1'b1;
in[159] : out[159] = 1'b1;
in[160] : out[160] = 1'b1;
in[161] : out[161] = 1'b1;
in[162] : out[162] = 1'b1;
in[163] : out[163] = 1'b1;
in[164] : out[164] = 1'b1;
in[165] : out[165] = 1'b1;
in[166] : out[166] = 1'b1;
in[167] : out[167] = 1'b1;
in[168] : out[168] = 1'b1;
in[169] : out[169] = 1'b1;
in[170] : out[170] = 1'b1;
in[171] : out[171] = 1'b1;
in[172] : out[172] = 1'b1;
in[173] : out[173] = 1'b1;
in[174] : out[174] = 1'b1;
in[175] : out[175] = 1'b1;
in[176] : out[176] = 1'b1;
in[177] : out[177] = 1'b1;
in[178] : out[178] = 1'b1;
in[179] : out[179] = 1'b1;
in[180] : out[180] = 1'b1;
in[181] : out[181] = 1'b1;
in[182] : out[182] = 1'b1;
in[183] : out[183] = 1'b1;
in[184] : out[184] = 1'b1;
in[185] : out[185] = 1'b1;
in[186] : out[186] = 1'b1;
in[187] : out[187] = 1'b1;
in[188] : out[188] = 1'b1;
in[189] : out[189] = 1'b1;
in[190] : out[190] = 1'b1;
in[191] : out[191] = 1'b1;
in[192] : out[192] = 1'b1;
in[193] : out[193] = 1'b1;
in[194] : out[194] = 1'b1;
in[195] : out[195] = 1'b1;
in[196] : out[196] = 1'b1;
in[197] : out[197] = 1'b1;
in[198] : out[198] = 1'b1;
in[199] : out[199] = 1'b1;
in[200] : out[200] = 1'b1;
in[201] : out[201] = 1'b1;
in[202] : out[202] = 1'b1;
in[203] : out[203] = 1'b1;
in[204] : out[204] = 1'b1;
in[205] : out[205] = 1'b1;
in[206] : out[206] = 1'b1;
in[207] : out[207] = 1'b1;
in[208] : out[208] = 1'b1;
in[209] : out[209] = 1'b1;
in[210] : out[210] = 1'b1;
in[211] : out[211] = 1'b1;
in[212] : out[212] = 1'b1;
in[213] : out[213] = 1'b1;
in[214] : out[214] = 1'b1;
in[215] : out[215] = 1'b1;
in[216] : out[216] = 1'b1;
in[217] : out[217] = 1'b1;
in[218] : out[218] = 1'b1;
in[219] : out[219] = 1'b1;
in[220] : out[220] = 1'b1;
in[221] : out[221] = 1'b1;
in[222] : out[222] = 1'b1;
in[223] : out[223] = 1'b1;
in[224] : out[224] = 1'b1;
in[225] : out[225] = 1'b1;
in[226] : out[226] = 1'b1;
in[227] : out[227] = 1'b1;
in[228] : out[228] = 1'b1;
in[229] : out[229] = 1'b1;
in[230] : out[230] = 1'b1;
in[231] : out[231] = 1'b1;
in[232] : out[232] = 1'b1;
in[233] : out[233] = 1'b1;
in[234] : out[234] = 1'b1;
in[235] : out[235] = 1'b1;
in[236] : out[236] = 1'b1;
in[237] : out[237] = 1'b1;
in[238] : out[238] = 1'b1;
in[239] : out[239] = 1'b1;
in[240] : out[240] = 1'b1;
in[241] : out[241] = 1'b1;
in[242] : out[242] = 1'b1;
in[243] : out[243] = 1'b1;
in[244] : out[244] = 1'b1;
in[245] : out[245] = 1'b1;
in[246] : out[246] = 1'b1;
in[247] : out[247] = 1'b1;
in[248] : out[248] = 1'b1;
in[249] : out[249] = 1'b1;
in[250] : out[250] = 1'b1;
in[251] : out[251] = 1'b1;
in[252] : out[252] = 1'b1;
in[253] : out[253] = 1'b1;
in[254] : out[254] = 1'b1;
in[255] : out[255] = 1'b1;
endcase
